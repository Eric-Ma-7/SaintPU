/* This is the ID stage of St.PU */
/*  */
`define InstOpBus 5:0
`define InstFuncBus 5:0
`define InstShamtBus 4:0
`define ImmBus 15:0
`define Enable 1'b1
`define Disable 1'b0

module ID(
input reg [`RegBus] pc_i,
input reg [`RegBus] inst_i,
input wire [`RegBus] reg1_data_i,
input wire [`RegBus] reg2_data_i,
/* Reset Signal */
input wire rst,
/* Ex data input enable */
input wire ex_wreg_i;
/* Ex data input destination addr */
input wire [`RegAddrBus] ex_wd_i;
/* EX data input*/
input wire [`RegBus] ex_wdata_i
/* Output Ports */
/* ALU Operation Code */
output reg [`AluOpBus] aluop_o,
/* ALU Opaeration Type Select */
output reg [`AluSelBus] alusel_o,
output reg [`RegBus] reg1_o,
output reg [`RegBus] reg2_o,
/* Write Destination */
output reg [`RegAddrBus] wd_o,
/* Write Enable */
output wire wreg_o,
/* Register Files Address */
output reg [`RegAddrBus] reg1_addr_o,
output reg [`RegAddrBus] reg2_addr_o,
/* Register Read Enable */
output wire reg1_read_o,
output wire reg2_read_o,
);
/* Internal Signals Define */
wire [`ImmBus] imm = inst_i[15:0];
wire [`InstOpBus] inst_op = inst_i[31:26];
wire [`InstFuncBus] inst_func = inst_i[5:0];
wire [`InstShamtBus] inst_sa = inst_i[10:6];
wire [`RegAddrBus] rs_addr = inst_i[25:21];
wire [`RegAddrBus] rt_addr = inst_i[20:16];
wire [`RegAddrBus] rd_addr = inst_i[15:11];
wire [`RegBus] sign_imm = {16{imm[15]},imm};
wire [`RegBus] unsign_imm = {16'h0,imm};
reg [`RegBus] imm_o;

always @(*) begin
    if (rst == `RstEnable) begin
        aluop_o = `EXE_NOP_OP;
        alusel_o = `EXE_RES_NOP;
        wd_o = `NOPRegAddr;
        wreg_o = `WriteDisable;
        reg1_read_o = `Disable;
        reg2_read_o = `Disable;
        reg1_addr_o = `NOPRegAddr;
        reg2_addr_o = `NOPRegAddr;
        imm_o = `ZeroWord;
    end else begin
        aluop_o = `EXE_NOP_OP;
        alusel_o = `EXE_RES_NOP;
        wd_o = rd_addr;
        reg1_read_o = `Disable;
        reg2_read_o = `Disable;
        reg1_addr_o = rs_addr;
        reg2_addr_o = rt_addr;
        imm_o = `ZeroWord;
        case (inst_op)
            `EXE_SPECIAL_INST:  begin
                case (inst_func)
                    `EXE_OR: begin
                        wreg_o = `WriteEnable;
                        aluop_o = `EXE_OR_OP;
                        alusel_o = ``EXE_RES_LOGIC;
                        reg1_read_o = `Enable;
                        reg2_read_o = `Enable;
                    end
                    `EXE_AND: begin
                        wreg_o = `WriteEnable;
                        aluop_o = `EXE_AND_OP;
                        alusel_o = `EXE_RES_LOGIC;
                        reg1_read_o = `Enable;
                        reg2_read_o = `Enable;
                    end
                    `EXE_XOR: begin
                        wreg_o = `WriteEnable;
                        aluop_o = `EXE_XOR_OP;
                        alusel_o = `EXE_RES_LOGIC;
                        reg1_read_o = `Enable;
                        reg2_read_o = `Enable;
                    end
                    `EXE_NOR: begin
                        wreg_o = `WriteEnable;
                        aluop_o = `EXE_NOR_OP;
                        alusel_o = `EXE_RES_LOGIC;
                        reg1_read_o = `Enable;
                        reg2_read_o = `Enable;
                    end
                    `EXE_SLLV: begin
                        wreg_o = `WriteEnable;
                        aluop_o = `EXE_SLL_OP;
                        alusel_o = `EXE_RES_SHIFT;
                        reg1_read_o = `Enable;
                        reg2_read_o = `Enable;
                    end
                    `EXE_SRLV: begin
                        wreg_o = `WriteEnable;
                        aluop_o = `EXE_SRL_OP;
                        alusel_o = `EXE_RES_SHIFT;
                        reg1_read_o = `Enable;
                        reg2_read_o = `Enable;
                    end
                    `EXE_SRAV: begin
                         wreg_o = `WriteEnable;
                        aluop_o = `EXE_SRA_OP;
                        alusel_o = `EXE_RES_SHIFT;
                        reg1_read_o = `Enable;
                        reg2_read_o = `Enable;
                    end
                    
                    default: begin
                    end
                endcase
                if (rs_addr == 5'h0) begin 
                    case (inst_func):
                        `EXE_SLL: begin
                            wreg_o = `WriteEnable;
                            aluop_o = `EXE_SLL_OP;
                            alusel_o = `EXE_RES_SHIFT;
                            reg1_read_o = `Disable;
                            reg2_read_o = `Enable;
                            imm_o = {27'h0,inst_sa};
                            wd_o = rd_addr;
                        end
                        `EXE_SRL: begin
                            wreg_o = `WriteEnable;
                            aluop_o = `EXE_SRL_OP;
                            alusel_o = `EXE_RES_SHIFT;
                            reg1_read_o = `Disable;
                            reg2_read_o = `Enable;
                            imm_o = {27'h0,inst_sa};
                            wd_o = rd_addr;
                        end
                        `EXE_SRA: begin
                            wreg_o = `WriteEnable;
                            aluop_o = `EXE_SRA_OP;
                            alusel_o = `EXE_RES_SHIFT;
                            reg1_read_o = `Disable;
                            reg2_read_o = `Enable;
                            imm_o = {27'h0,inst_sa};
                            wd_o = rd_addr;
                        end
                    endcase
                end
            end
            `EXE_ORI: begin
                wreg_o = `WriteEnable;
                aluop_o = `EXE_OR_OP;
                alusel_o = `EXE_RES_LOGIC;
                reg1_read_o = `Enable;
                reg2_read_o = `Disable;
                imm_o = unsign_imm;
                wd_o =  rt_addr;
            end
            `EXE_ANDI: begin
                wreg_o = `WriteEnable;
                aluop_o = `EXE_AND_OP;
                alusel_o = `EXE_RES_LOGIC;
                reg1_read_o = `Enable;
                reg2_read_o = `Disable;
                imm_o = unsign_imm;
                wd_o =  rt_addr;
            end
            `EXE_XORI: begin
                wreg_o = `WriteEnable;
                aluop_o = `EXE_XOR_OP;
                alusel_o = `EXE_RES_LOGIC;
                reg1_read_o = `Enable;
                reg2_read_o = `Disable;
                imm_o = unsign_imm;
                wd_o =  rt_addr;
            end
            `EXE_LUI: begin
                wreg_o = `WriteEnable;
                aluop_o = `EXE_OR_OP;
                alusel_o = `EXE_RES_LOGIC;
                reg1_read_o = `Disable;
                reg2_read_o = `Disable;
                imm_o = {imm,16'h0};
                wd_o = rt_addr;
            end
            
            default: begin
            end
        endcase
end

always @(*) begin
    if (rst == `RstEnable) begin
        reg1_o =  `ZeroWord;
    end else if ((ex_wreg_i == `Enable) && (ex_wd_i == reg1_addr_o) && (reg1_read_o == `Enable)) begin
        reg1_o = ex_wdata_i;
    end else if ((reg1_read_o == `Enable) && (mem_wreg_i == `Enable) && (mem_wd_i == reg1_addr_o
    )) begin
        reg1_o = mem_wdata_i;
    end else if (reg1_read_o == `Enable) begin
        reg1_o = reg1_data_i;
    end else if (reg1_read_o == `Disable) begin
        reg1_o = imm_o;
    end else begin
        reg1_o = `ZeroWord;
    end
end

always @(*) begin
    if (rst == `RstEnable) begin
        reg2_o =  `ZeroWord;
    end else if ((ex_wreg_i == `Enable) && (ex_wd_i == reg1_addr_o) && (reg2_read_o == `Enable)) begin
        reg2_o = ex_wdata_i;
    end else if ((reg2_read_o == `Enable) && (mem_wreg_i == `Enable) && (mem_wd_i == reg2_addr_o
    )) begin
        reg2_o = mem_wdata_i;
    end else if (reg1_read_o == `Enable) begin
        reg2_o = reg1_data_i;
    end else if (reg1_read_o == `Disable) begin
        reg2_o = imm_o;
    end else begin
        reg2_o = `ZeroWord;
    end
end

endmodule